--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:    23:28:04 07/14/05
-- Design Name:    
-- Module Name:    set_rgb - Behavioral
-- Project Name:   
-- Target Device:  
-- Tool versions:  
-- Description:
--
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
--------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

---- Uncomment the following library declaration if instantiating
---- any Xilinx primitives in this chiffre.
--library UNISIM;
--use UNISIM.VComponents.all;

-- ************************************************
-- ******************** ENTITE ********************
-- ************************************************

entity set_rgb is
	PORT(
			Clk : in std_logic;
-- Ports qui renvoient les coordonns du pointeur
			X : IN std_logic_vector(9 downto 0);
			Y : IN std_logic_vector(9 downto 0);
-- Port qui permet de savoir si l'on se situe dans la zone d'affichage ou non
			VIDEO_EN : IN std_logic	;
-- Ports l'acquisition des joysticks
			red_btn : IN std_logic;
			green_btn : IN std_logic;
			yellow_btn : IN std_logic;
			blue_btn : IN std_logic;
			game_over  : IN std_logic;
-- Ports concernent le mouvenent de la balle et des raquettes
			--CLK_Ball : IN std_logic;
			--CLK_raquette : IN std_logic;
			
			
--PAUSE_ENABLED : IN std_logic;
-- Ports sur lesquels, on dfinie la couleur du pixel  afficher
 			R : out std_logic;
      	G : out std_logic;
      	B : out std_logic
		 );

end set_rgb;  

-- ******************************************************
-- ******************** ARCHITECTURE ********************
-- ******************************************************

architecture Hamid of set_rgb is

---------------------------------------------------------			  								  								  								 
--------- DECLARATION DES SIGNAUX ET CONSTANTES ---------
---------------------------------------------------------

																																	   
--	DEFINTION DES CONSTANTES 0,1,2,3,4,5,6,7,8,9 UTILISANT LE TABLEAU "CHIFFRE"
------------------------------------------------------------------------------

	type chiffre is array (0 to 39, 0 to 19) of natural; 

	constant zero: chiffre:=		((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));
							  	
	constant un: chiffre:=			((0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0),
  											(0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0));

	constant deux: chiffre:=		((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));

 	constant	trois: chiffre:=		((0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),	
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
						   				(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));


  constant quatre: chiffre:=		((1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1));


	constant	cinq: chiffre:=		((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));

	constant	six: chiffre:=			((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));
										

	constant	sept: chiffre:=		((1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0));
			  	
	constant	huit: chiffre:=		((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
 											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
 											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));
										
									
	constant	neuf: chiffre:=		((0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
 											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0),
											(0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0),
 											(1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0));


-- DEFINITION D'UN TABLEAU (40,70) POUR AFFICHER "WIN"
------------------------------------------------------

	type wini is array (0 to 39, 0 to 69) of natural;			 

  	constant win: wini:=				((1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1),
											(0,0,0,1,0,0,0,0,0,1,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1),
											(0,0,0,1,0,0,0,0,1,0,0,1,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1),
											(0,0,0,0,1,0,0,1,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1),
											(0,0,0,0,1,0,1,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1),
 											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1));
		  	
-- DEFINITION D'UN TABLEAU (40,110) POUR AFFICHER "LOSE"
--------------------------------------------------------

	type losed is array (0 to 39, 0 to 109) of natural;

	constant lose: losed:=			((1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
 											(0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));
			  	






	type debu2 is array (0 to 39, 0 to 179) of natural;
  	constant debu: debu2  :=   	((1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
 											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0),
 											(0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1,1));






	type restart is array (0 to 19, 0 to 157) of natural;

	constant start: restart:=		((1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1),
 											(1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1),
											(1,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0),
											(1,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,1,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,0,0,1,0,0,0,0),
											(1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,0,0,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0),
 											(1,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,1,1,0,0,0,0,0,0,0,1,1,1,1,1,1,1,1,1,1,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,0,0));


-- DEFINITION D'UN TABLEAU (5,15) POUR AFFICHER LE MISSILE
----------------------------------------------------------

	type miss is array (0 to 4, 0 to 14) of natural;

-- LANCE PAR LE JOUEUR A

	constant missile_A: miss:=		((1,1,1,1,1,1,1,1,1,0,0,0,0,0,0),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(0,0,0,0,0,0,0,1,1,1,1,1,1,1,1),
											(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
											(1,1,1,1,1,1,1,1,1,0,0,0,0,0,0));
-- LANCE PAR LE JOUEUR B
				  	
	constant missile_B: miss:=		((0,0,0,0,0,0,1,1,1,1,1,1,1,1,1),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(1,1,1,1,1,1,1,1,0,0,0,0,0,0,0),
											(0,0,0,0,0,1,0,0,0,0,0,0,0,0,0),
											(0,0,0,0,0,0,1,1,1,1,1,1,1,1,1));
												  
-- DEFINITION D'UN TABLEAU (15,15) POUR AFFICHER L'EXPLOSION DU MISSILE
-----------------------------------------------------------------------

	type explo is array (0 to 14, 0 to 14) of natural;

-- SUR LE JOUEUR A
	
	constant explose_A: explo:=	((1,1,1,0,0,0,0,0,0,0,0,0,0,0,0),
											(0,0,0,1,1,0,0,0,0,0,0,0,0,0,0),
  										   (0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
  									    	(0,0,0,0,0,0,0,0,0,1,0,0,0,0,0),
  									    	(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  									   	(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  								   	   (0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
  									      (0,0,0,0,0,1,1,0,0,0,0,0,0,0,0),
  									    	(0,0,0,1,1,0,0,0,0,0,0,0,0,0,0), 
  									      (1,1,1,0,0,0,0,0,0,0,0,0,0,0,0));
-- SUR LE JOUEUR B  									    

	constant explose_B: explo:= 	((0,0,0,0,0,0,0,0,0,0,0,0,0,1,1),
  										   (0,0,0,0,0,0,0,0,0,0,0,1,1,0,0),
  										   (0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
  										   (0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
  										   (0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
  									    	(0,0,0,0,0,0,1,0,0,0,0,0,0,0,0),
  									    	(0,0,0,0,0,0,0,1,0,0,0,0,0,0,0),
  									   	(0,0,0,0,0,0,0,0,1,0,0,0,0,0,0),
  								   	   (0,0,0,0,0,0,0,0,0,1,1,0,0,0,0),
  									      (0,0,0,0,0,0,0,0,0,0,1,0,0,0,0),
  									    	(0,0,0,0,0,0,0,0,0,0,0,1,1,0,0), 
  									      (0,0,0,0,0,0,0,0,0,0,0,0,0,1,1));
  									    
-- *********************************************************************************************************

    
-- COORDONNEES DU POINTEUR DE TYPE ENTIER

	signal iX,iY : integer range 0 to 1023;	
 	-- Variables du chronomtres
	--changed
	signal second_lower_digit: integer range 0 to 10 := 9;
	signal second_upper_digit: integer range 0 to 10 := 5;
	signal minutes: integer range 0 to 10 := 3;
	signal cpt: integer range 0 to 10000000 := 0;		
   signal miliseconds : integer range 0 to 10 := 9;

-- COORDONNEES Y DES RAQUETTES

	signal y_raquette_A,y_raquette_B: integer range 0 to 1023:=200; 

-- CONTROLE DE LA BALLE

	signal xb,yb : integer range 0 to 1023;		  						 -- Coordonnes (x,y) de la balle
	signal dirX,dirY: std_logic;						   					 -- Dtermine sa direction
   -- AFFICHAGE ET COORDONNEES DU CHAMPIGNION
	signal clk_champignion: std_logic_vector(19 downto 0);
	signal x_champignion: integer range 0 to 1023 := 200;
	signal y_champignion: integer range 0 to 1023 := 200;
	signal champignion_affiche: std_logic := '1';
	-- GARDER TRACE DU DRENIERE RAQUETTE QUI A FRAPPE LA BALLE
	type JOUEUR is (JOUEUR_A, JOUEUR_B);
	signal raquette_source: JOUEUR;
	signal clk_creation_champignion : std_logic_vector(19 downto 0):= "00000000000000000000";
-- CONTROLE DES SCORES ET DE LA FIN DE LA PARTIE

	signal score_A,score_B : integer range 0 to 1023:= 0;				 -- Score du joueur A et du joueur B
	signal x_lose, x_win: integer range 0 to 1023;						 -- variable de positionnement du "gagant" et du "perdant" de la partie

-- DEFINTIION DES SIGNAUX NECESSAIRES AU CONTROLE DES MISSILES

	signal x_missile_A: integer range 0 to 1023:=20;					 -- |
	signal y_missile_A: integer range 0 to 1023:=10;	 				 -- |	Coordonnes des missiles lancs par
	signal x_missile_B: integer range -20 to 1023:=605;				 -- |	le joueur A et le joueur B
	signal y_missile_B: integer range 0 to 1023:=10;					 -- |
						 
 	signal missileA_enable, missileB_enable: std_logic:='0';			 
	signal explosion_A, explosion_B: std_logic:='0';
																				
-- DEFINITION DE LA PALETTE DES 8 COULEURS POUR L'AFFICHAGE

	signal pixel_enable: std_logic;
	signal pixel_white: std_logic;								  
	signal pixel_yellow: std_logic;
	signal pixel_blue: std_logic;
	signal pixel_green: std_logic;																					  
	signal pixel_red: std_logic;
	signal pixel_cyan: std_logic;
	signal pixel_magenta: std_logic;

-- DEFINITION DE L'ETAT DE LA PARTIE

	type PARTIE is (DEBUT,EN_COURS,FIN,PAUSE);
	signal ETAT_PARTIE : PARTIE;

	signal yy: integer range 0 to 1023:=600;
   
	
-- *******************************************************************************************************
-- *******************************************************************************************************
-- ***************************************** DEBUT DU PROGRAMME ******************************************
-- *******************************************************************************************************
-- *******************************************************************************************************

begin								
																			
	iX<=CONV_INTEGER(X);		-- conversion des coordonnes binaires (X,Y) du pointeur en ENTIER									 
	iY<=CONV_INTEGER(Y);

-- *******************************************************************************************************
-- ******** DEPLACEMENT DES RAQUETTES, CONTROLE DE L'ETAT DES MISSILES ET DE L'ETAT DE LA PARTIE *********
-- *******************************************************************************************************


------------------------------------------------------------------------------										 
---------- CONTROLE DE L'ETAT DE LA PARTIE : DEBUT, EN COURS ET FIN ----------
------------------------------------------------------------------------------	
	
	
	CTRL_CHRONO: process(CLK)
	begin
		if CLK'event and CLK='1' then
			if ETAT_PARTIE = DEBUT then
				miliseconds <= 9;
				second_lower_digit <= 9;
				second_upper_digit <= 5;
				minutes <= 3;
			end if;
			if ETAT_PARTIE = EN_COURS then
				cpt <=cpt+1;
				if cpt = 10000000 then
					cpt <= 0;
					miliseconds <= miliseconds - 1;
					--if miliseconds = 0 then
						miliseconds <= 9;
						second_lower_digit  <= second_lower_digit -1;
						if second_lower_digit = 0 then
							second_lower_digit <= 9;
							second_upper_digit <=  second_upper_digit -1;
							if second_upper_digit = 0 then
								second_upper_digit <= 5;
								minutes <= minutes -1 ;
							end if;
						end if;
					--end if;
					
				end if;
			end if;
		end if;
	end process;
 	

 	
-- ********************************************************************************************************
-- *************************** PROCESS DU MOUVEMENT DE LA BALLE ET DES MISSILES ***************************
-- ********************************************************************************************************
 
	

-- *******************************************************************************************************
-- *************** PROCESS SENSIBLE AU POINTEUR : AFFICHAGE D'UN PIXEL (iX,iY) SUR L'ECRAN ***************
-- *******************************************************************************************************

	DRAW_DISP : process(iX,iY,red_btn,green_btn,yellow_btn,blue_btn)
	begin

---------------------------------------------------------
---------- INITIALISATION DU COLOR PIXEL A '0' ----------
---------------------------------------------------------

		pixel_enable<='0';
		pixel_white<='0';
		pixel_cyan<='0';
		pixel_magenta<='0';
		pixel_yellow<='0';
		pixel_green<='0';
		pixel_blue<='0';
		pixel_red<='0';

----------------------------------------
---------- AFFICHAGE DES CARREAUX ----------
----------------------------------------
		
		if iX<310 and iX>10 and iY>10 and iY<230 then
		
			pixel_blue<='1';
			if blue_btn='1' then
				pixel_enable<='1';
			end if;
		
		end if;
		
	if iX<629 and iX>330 and iY>10 and iY<230 then
		
			pixel_green<='1';
			if green_btn='1' then
				pixel_enable<='1';
			end if;											
		
		end if;
		
		if iX<310 and iX>10 and iY>250 and iY<469 then
		
			pixel_red<='1';
			if red_btn='1' then
				pixel_enable<='1';
			end if;											
		
		end if;
		
		if iX<629 and iX>330 and iY>250 and iY<469 then
		
			pixel_yellow<='1';
			if yellow_btn='1' then
				pixel_enable<='1';
			end if;											
		
		end if;
---------------------------------------------------------------
---------- AFFICHAGE DU CADRE (LIMITES DE LA PARTIE) ----------
---------------------------------------------------------------

		if iX=0 or iX=639 or iY=0 or iY=479 then
 			pixel_enable<='1';
			pixel_blue<='1';
		end if;

---------------------------------------------------			  								  								  								 
--------- AFFICHAGE DE LA PHRASE: Lose ---------
---------------------------------------------------

		if game_over='1' and iY>219 and iY<261 and iX<374 and iX>264 and lose(iY-220, iX-265)=1 then
			pixel_red <= '1';
			pixel_enable <= '1';
		end if;

-----------------------------------------------------------------------------			  								  								  								 
--------- PALETTE VIDEO : ACTIVATION DU PIXEL DE COORDONNEE (iX,iY) ---------
-----------------------------------------------------------------------------
end process;

process(VIDEO_EN, pixel_enable, pixel_white, pixel_yellow,pixel_blue,pixel_green,pixel_red,pixel_cyan,pixel_magenta)
begin
		  if VIDEO_EN='1' and pixel_enable='1' then
		     
			  if pixel_white='1' then
			    R <='1'; G <='1'; B <='1';			-- BLANC
	   	  end if;
																				  
 			  if pixel_yellow='1' then					-- JAUNE
				 R <='1'; G <='1'; B <='0';
			  end if;

			  if pixel_blue='1' then					-- BLEU
			  	 R <='0'; G <='0'; B <='1';
			  end if;

			  if pixel_green='1' then					-- VERT
			  	 R <='0'; G <='1'; B <='0';
			  end if;			
			 													
			  if pixel_red='1' then						-- ROUGE
				 R <='1'; G <='0'; B <='0';
			  end if;

			  if pixel_cyan='1' then					-- CYAN
			  	 R <='0'; G <='1'; B <='1';
			  end if;

			  if pixel_magenta='1' then				-- MAGENTA
			  	 R <='1'; G <='0'; B <='1';
			  end if;

			 else
			 
			    R <='0'; G <='0'; B <='0';		   -- NOIR 
   		  
		  end if;							  
		
end process;

	
end Hamid;
																	